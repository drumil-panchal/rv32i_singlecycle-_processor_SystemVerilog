//------------------------------------------
//resgister file
//------------------------------------------

import risc_pkg::*;
module registerfile(
    input logic clk,
    input logic reset_n,
    
    input logic [4:0] rs1_addr,
    input logic [4:0] rs2_addr,
    input logic [4:0] rd_addr,
    
    input logic rf_wr_en,
    input logic [31:0] wr_data,
    
    output logic [31:0] rs1_data,
    output logic [31:0] rs2_data
    );
    
    logic [31:0] regs[0:31];                    //register file of 32x32
    integer i;
    
    //read logic
    assign rs1_data = regs[rs1_addr];
    assign rs2_data = regs[rs2_addr];
    
    //write logic
    always_ff @(posedge clk or negedge reset_n) begin  
    
        if(!reset_n) begin
            for(i=0; i<32; i++)
                regs[i] <= 32'd0;                                                      //reset all registers to 0
        end
        
        else if (rf_wr_en && (rd_addr != 5'd0)) begin                  //if write enable is high and destination address is not 0
            regs[rd_addr] <= wr_data;
        end
    end 
    
endmodule
